
module boolean_functions (
input wire A,
input wire B,
input wire C,
input wire D,
output wire F
);
assign F = (~A & B) | (C & D) | (A & ~D);
endmodule